`define KNN_ADDR_W 3  //address width
`define KNN_WDATA_W 32 //write data width // ERIC: Changed to accomodate 32 bit words
`ifndef DATA_W
 `define DATA_W 32      //cpu data width
`endif
